module hexdisplay(

	output		     [7:0]		HEX,
	input				  [3:0]		I
);



//=======================================================
//  REG/WIRE declarations
//=======================================================

	


//=======================================================
//  Structural coding
//=======================================================

	assign HEX[0] = (~I[3]&I[2]&~I[1]&~I[0]) + (I[3]&~I[2]&I[1]&I[0]) + (I[3]&I[2]&~I[1]&I[0]);
	assign HEX[1] = (~I[3]&I[2]&~I[1]&I[0]) + (~I[3]&I[2]&I[1]&~I[0]) + (I[3]&~I[2]&I[1]&I[0]) + (I[3]&I[2]&~I[1]&~I[0]) + (I[3]&I[2]&I[1]&~I[0]) + (I[3]&I[2]&I[1]&I[0]);
	assign HEX[2] = (~I[3]&~I[2]&~I[1]&I[0]) + (~I[3]&~I[2]&I[1]&~I[0]) + (I[3]&I[2]&~I[1]&~I[0]) + (I[3]&I[2]&I[1]&~I[0]) + (I[3]&I[2]&I[1]&I[0]);
	assign HEX[3] = (~I[3]&~I[2]&~I[1]&I[0]) + (~I[3]&I[2]&~I[1]&~I[0]) + (~I[3]&I[2]&I[1]&I[0]) + (I[3]&~I[2]&I[1]&~I[0]) + (I[3]&I[2]&I[1]&I[0]);
	assign HEX[4] = (~I[3]&~I[2]&~I[1]&I[0]) + (~I[3]&~I[2]&I[1]&I[0]) + (~I[3]&I[2]&~I[1]&~I[0]) + (~I[3]&I[2]&~I[1]&I[0]) + (~I[3]&I[2]&I[1]&I[0]) + (I[3]&~I[2]&~I[1]&I[0]);
	assign HEX[5] = (~I[3]&~I[2]&~I[1]&I[0]) + (~I[3]&~I[2]&I[1]&~I[0]) + (~I[3]&~I[2]&I[1]&I[0]) + (~I[3]&I[2]&I[1]&I[0]) + (I[3]&I[2]&~I[1]&I[0]);
	assign HEX[6] = (~I[3]&~I[2]&~I[1]&~I[0]) + (~I[3]&~I[2]&~I[1]&I[0]) + (~I[3]&I[2]&I[1]&I[0]) + (I[3]&I[2]&~I[1]&~I[0]);
		
	
endmodule
